`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/27/2025 10:46:45 AM
// Design Name: 
// Module Name: cricketGame
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////




module cricketGame(
    input clk_fpga,
    input reset,
    input play,
    input teamSwitch,
    output [7:0] binaryruns,
    output [3:0] binarywickets,
    output [15:0] leds,
    output inningOver,
    output gameOver,
    output winner
);

    // Internal wires
    wire [11:0] team1Data;      // stores and updates team1's runs and wickets when switch is 0
    wire [11:0] team2Data;      // stores and updates team2's runs and wickets when switch is 1
    wire [6:0] team1Balls;      // number of team1's deliveries that are legal balls, shown on LEDs
    wire [6:0] team2Balls;      // number of team2's deliveries that are legal balls, shown on LEDs
    wire [3:0] lfsr_out;        // pseudo-random number from linear feedback shift register

    // Pseudo random number generator using a linear feedback shift register
    lfsr1 g1(clk_fpga, reset, lfsr_out); // 4-bit LFSR output used as a signal/event generator

    // Assign scores and wickets based on pseudo random number generated by lfsr
    score_and_wickets g2(
        clk_fpga, reset, play, teamSwitch, lfsr_out,
        gameOver, binaryruns, binarywickets, team1Data, team2Data
    );

    // Comparator that finds and locks in the winner when the game is over
    score_comparator g3(
        clk_fpga, reset, team1Data, team2Data, team1Balls, team2Balls,
        binarywickets, leds, inningOver, gameOver, winner
    );

    // Assign LEDs based on balls of team in play, or scrolls winner when game is over
    led_controller g4(
        clk_fpga, reset, teamSwitch, play, lfsr_out,
        inningOver, gameOver, leds, team1Balls, team2Balls
    );

endmodule





